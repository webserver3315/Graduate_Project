module my_and
		(
		input a, b,
		output c
		);
	assign c = a&b;
endmodule
