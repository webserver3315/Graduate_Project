// DESCRIPTION: Verilator: Verilog example module
//
// This file ONLY is placed under the Creative Commons Public Domain, for
// any use, without warranty, 2017 by Wilson Snyder.
// SPDX-License-Identifier: CC0-1.0

// See also https://verilator.org/guide/latest/examples.html"
`include "Black_Cell.v"

module top
   (
      input clk
   );
   initial begin
      $display("Hello World!");
      $finish;
   end
endmodule
